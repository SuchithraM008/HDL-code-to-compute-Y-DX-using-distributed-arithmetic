module ROM(S,Count,Y);

input [7:0]S;
input [4:0] Count;
output [10:0]Y;
reg [9:0]R[15:0][15:0];

// ROM1
assign R[0][0]=10'd0;
assign R[1][0]=10'd45;
assign R[2][0]=10'd45;
assign R[3][0]=10'd90;
assign R[4][0]=10'd45;
assign R[5][0]=10'd90;
assign R[6][0]=10'd90;
assign R[7][0]=10'd135;
assign R[8][0]=10'd45;
assign R[9][0]=10'd90;
assign R[10][0]=10'd90;
assign R[11][0]=10'd135;
assign R[12][0]=10'd90;
assign R[13][0]=10'd135;
assign R[14][0]=10'd135;
assign R[15][0]=10'd180;

//ROM2
assign R[0][1]=10'd0;
assign R[1][1]=10'd45;
assign R[2][1]=10'd45;
assign R[3][1]=10'd90;
assign R[4][1]=10'd45;
assign R[5][1]=10'd90;
assign R[6][1]=10'd90;
assign R[7][1]=10'd135;
assign R[8][1]=10'd45;
assign R[9][1]=10'd90;
assign R[10][1]=10'd90;
assign R[11][1]=10'd135;
assign R[12][1]=10'd90;
assign R[13][1]=10'd135;
assign R[14][1]=10'd135;
assign R[15][1]=10'd180;

// ROM3
assign R[0][2]=10'd0;
assign R[1][2]=10'd63;
assign R[2][2]=10'd53;
assign R[3][2]=10'd116;
assign R[4][2]=10'd36;
assign R[5][2]=10'd99;
assign R[6][2]=10'd89;
assign R[7][2]=10'd152;
assign R[8][2]=10'd12;
assign R[9][2]=10'd75;
assign R[10][2]=10'd65;
assign R[11][2]=10'd128;
assign R[12][2]=10'd48;
assign R[13][2]=10'd111;
assign R[14][2]=10'd101;
assign R[15][2]=10'd164;

// ROM4
assign R[0][3]=-10'd0;
assign R[1][3]=-10'd12;
assign R[2][3]=-10'd36;
assign R[3][3]=-10'd48;
assign R[4][3]=-10'd53;
assign R[5][3]=-10'd65;
assign R[6][3]=-10'd89;
assign R[7][3]=-10'd101;
assign R[8][3]=-10'd63;
assign R[9][3]=-10'd75;
assign R[10][3]=-10'd99;
assign R[11][3]=-10'd111;
assign R[12][3]=-10'd116;
assign R[13][3]=-10'd128;
assign R[14][3]=-10'd152;
assign R[15][3]=-10'd164;

//ROM5
assign R[0][4]=10'd0;
assign R[1][4]=10'd59;
assign R[2][4]=10'd24;
assign R[3][4]=10'd83;
assign R[4][4]=-10'd24;
assign R[5][4]=10'd35;
assign R[6][4]=10'd0;
assign R[7][4]=10'd59;
assign R[8][4]=-10'd59;
assign R[9][4]=10'd0;
assign R[10][4]=-10'd35;
assign R[11][4]=10'd24;
assign R[12][4]=-10'd83;
assign R[13][4]=-10'd24;
assign R[14][4]=-10'd59;
assign R[15][4]=10'd0;

// ROM6
assign R[0][5]=10'd0;
assign R[1][5]=-10'd59;
assign R[2][5]=-10'd24;
assign R[3][5]=-10'd83;
assign R[4][5]=10'd24;
assign R[5][5]=-10'd35;
assign R[6][5]=10'd0;
assign R[7][5]=-10'd59;
assign R[8][5]=10'd59;
assign R[9][5]=10'd0;
assign R[10][5]=10'd35;
assign R[11][5]=-10'd24;
assign R[12][5]=10'd83;
assign R[13][5]=10'd24;
assign R[14][5]=10'd59;
assign R[15][5]=10'd0;

// ROM7
assign R[0][6]=10'd0;
assign R[1][6]=10'd53;
assign R[2][6]=-10'd12;
assign R[3][6]=10'd41;
assign R[4][6]=-10'd63;
assign R[5][6]=-10'd10;
assign R[6][6]=-10'd75;
assign R[7][6]=-10'd22;
assign R[8][6]=-10'd36;
assign R[9][6]=10'd17;
assign R[10][6]=-10'd48;
assign R[11][6]=10'd5;
assign R[12][6]=-10'd99;
assign R[13][6]=-10'd46;
assign R[14][6]=-10'd111;
assign R[15][6]=-10'd58;

//ROM8
assign R[0][7]=10'd0;
assign R[1][7]=10'd36;
assign R[2][7]=10'd63;
assign R[3][7]=10'd99;
assign R[4][7]=10'd12;
assign R[5][7]=10'd48;
assign R[6][7]=10'd75;
assign R[7][7]=10'd111;
assign R[8][7]=-10'd53;
assign R[9][7]=-10'd17;
assign R[10][7]=10'd10;
assign R[11][7]=10'd46;
assign R[12][7]=-10'd41;
assign R[13][7]=-10'd5;
assign R[14][7]=10'd22;
assign R[15][7]=10'd58;

// ROM9
assign R[0][8]=10'd0;
assign R[1][8]=10'd45;
assign R[2][8]=-10'd45;
assign R[3][8]=10'd0;
assign R[4][8]=-10'd45;
assign R[5][8]=10'd0;
assign R[6][8]=-10'd90;
assign R[7][8]=-10'd45;
assign R[8][8]=10'd45;
assign R[9][8]=10'd90;
assign R[10][8]=10'd0;
assign R[11][8]=10'd45;
assign R[12][8]=10'd0;
assign R[13][8]=10'd45;
assign R[14][8]=-10'd45;
assign R[15][8]=10'd0;

// ROM10
assign R[0][9]=10'd0;
assign R[1][9]=10'd45;
assign R[2][9]=-10'd45;
assign R[3][9]=10'd0;
assign R[4][9]=-10'd45;
assign R[5][9]=10'd0;
assign R[6][9]=-10'd90;
assign R[7][9]=-10'd45;
assign R[8][9]=10'd45;
assign R[9][9]=10'd90;
assign R[10][9]=10'd0;
assign R[11][9]=10'd45;
assign R[12][9]=10'd0;
assign R[13][9]=10'd45;
assign R[14][9]=-10'd45;
assign R[15][9]=10'd0;

// ROM11
assign R[0][10]=10'd0;
assign R[1][10]=10'd36;
assign R[2][10]=-10'd63;
assign R[3][10]=-10'd27;
assign R[4][10]=10'd12;
assign R[5][10]=10'd48;
assign R[6][10]=-10'd51;
assign R[7][10]=-10'd15;
assign R[8][10]=10'd53;
assign R[9][10]=10'd89;
assign R[10][10]=-10'd10;
assign R[11][10]=10'd26;
assign R[12][10]=10'd65;
assign R[13][10]=10'd101;
assign R[14][10]=10'd2;
assign R[15][10]=10'd38;

// ROM12
assign R[0][11]=10'd0;
assign R[1][11]=-10'd53;
assign R[2][11]=-10'd12;
assign R[3][11]=-10'd65;
assign R[4][11]=10'd63;
assign R[5][11]=10'd10;
assign R[6][11]=10'd51;
assign R[7][11]=-10'd2;
assign R[8][11]=-10'd36;
assign R[9][11]=-10'd89;
assign R[10][11]=-10'd48;
assign R[11][11]=-10'd101;
assign R[12][11]=10'd27;
assign R[13][11]=-10'd26;
assign R[14][11]=10'd15;
assign R[15][11]=-10'd38;

// ROM13
assign R[0][12]=10'd0;
assign R[1][12]=10'd24;
assign R[2][12]=-10'd59;
assign R[3][12]=-10'd35;
assign R[4][12]=10'd59;
assign R[5][12]=10'd83;
assign R[6][12]=10'd0;
assign R[7][12]=10'd24;
assign R[8][12]=-10'd24;
assign R[9][12]=10'd0;
assign R[10][12]=-10'd83;
assign R[11][12]=-10'd59;
assign R[12][12]=10'd35;
assign R[13][12]=10'd59;
assign R[14][12]=-10'd24;
assign R[15][12]=10'd0;

// ROM14
assign R[0][13]=-10'd0;
assign R[1][13]=-10'd24;
assign R[2][13]=10'd59;
assign R[3][13]=10'd35;
assign R[4][13]=-10'd59;
assign R[5][13]=-10'd83;
assign R[6][13]=-10'd0;
assign R[7][13]=-10'd24;
assign R[8][13]=10'd24;
assign R[9][13]=-10'd0;
assign R[10][13]=10'd83;
assign R[11][13]=10'd59;
assign R[12][13]=-10'd35;
assign R[13][13]=-10'd59;
assign R[14][13]=10'd24;
assign R[15][13]=-10'd0;

// ROM15
assign R[0][14]=10'd0;
assign R[1][14]=10'd12;
assign R[2][14]=-10'd36;
assign R[3][14]=-10'd24;
assign R[4][14]=10'd53;
assign R[5][14]=10'd65;
assign R[6][14]=10'd17;
assign R[7][14]=10'd29;
assign R[8][14]=-10'd63;
assign R[9][14]=-10'd51;
assign R[10][14]=-10'd99;
assign R[11][14]=-10'd87;
assign R[12][14]=-10'd10;
assign R[13][14]=10'd2;
assign R[14][14]=-10'd46;
assign R[15][14]=-10'd34;

// ROM16
assign R[0][15]=10'd0;
assign R[1][15]=10'd63;
assign R[2][15]=-10'd53;
assign R[3][15]=10'd10;
assign R[4][15]=10'd36;
assign R[5][15]=10'd99;
assign R[6][15]=-10'd17;
assign R[7][15]=10'd46;
assign R[8][15]=-10'd12;
assign R[9][15]=10'd51;
assign R[10][15]=-10'd65;
assign R[11][15]=-10'd2;
assign R[12][15]=10'd24;
assign R[13][15]=10'd87;
assign R[14][15]=-10'd29;
assign R[15][15]=10'd34;

Add_Sub_Nbit #(.N(10)) Call_1 (.A(R[(S[3:0])][Count+Count]),.B(R[(S[7:4])][Count+Count+1'b1]),.k(1'b0),.S(Y));


endmodule
